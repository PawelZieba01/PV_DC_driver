PWM RC filter 2

VSUPPLY VCC 0 5V
C2 VCC 0 100n

X1 P_IN N_IN VCC 0 OUT LM324

VPWM VIN 0 PULSE 0 0.1 0 0 0 25u 50u

R3 VIN P_IN 1600
C3 P_IN 0 100n

R2 0 N_IN 410
R1 OUT N_IN 10k
C1 N_IN OUT 100n


.TRAN 0 5m 0 1u
.PROBE
.LIB "EVAL_TOS.LIB"
.END
